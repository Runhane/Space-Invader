module press_fire_text_map
(
	input logic [5:0] X,
	input logic [4:0] Y,
	output logic pixel
);

	logic [7:0] rom_address;
	logic [7:0] text_slice;
	
	assign pixel = text_slice[3'b111 - X[2:0]];
	
	press_fire_rom pfr(.address(rom_address), .data(text_slice));

	always_comb begin
	
		if(X >= 6'd0 && X < 6'd8 && Y >= 5'd0 && Y < 5'd16)
			rom_address = 8'd0 + Y;
		
		else if(X >= 6'd8 && X < 6'd16 && Y >= 5'd0 && Y < 5'd16)
			rom_address = 8'd16 + Y;
		
		else if(X >= 6'd16 && X < 6'd24 && Y >= 5'd0 && Y < 5'd16)
			rom_address = 8'd32 + Y;
		
		else if(X >= 6'd24 && X < 6'd32 && Y >= 5'd0 && Y < 5'd16)
			rom_address = 8'd48 + Y;
			
		else if(X >= 6'd32 && X < 6'd40 && Y >= 5'd0 && Y < 5'd16)
			rom_address = 8'd64 + Y;
			
		else if(X >= 6'd40 && X < 6'd48 && Y >= 5'd0 && Y < 5'd16)
			rom_address = 8'd80 + Y;
			
		else if(X >= 6'd48 && X < 6'd56 && Y >= 5'd0 && Y < 5'd16)
			rom_address = 8'd96 + Y;
			
		
		
		
		else if(X >= 6'd8 && X < 6'd16 && Y >= 5'd16)
			rom_address = 8'd128 + Y - 8'd16;
		
		else if(X >= 6'd16 && X < 6'd24 && Y >= 5'd16)
			rom_address = 8'd144 + Y - 8'd16;
	
		else if(X >= 6'd24 && X < 6'd32 && Y >= 5'd16)
			rom_address = 8'd160 + Y - 8'd16;
		
		else if(X >= 6'd32 && X < 6'd40 && Y >= 5'd16)
			rom_address = 8'd176 + Y - 8'd16;
		
		else if(X >= 6'd40 && X < 6'd48 && Y >= 5'd16)
			rom_address = 8'd192 + Y - 8'd16;
		else
			rom_address = 8'd176 + Y - 8'd16;	
		
	end

endmodule 

module press_fire_rom
(
	input [7:0] address,
	output [7:0] data
);

	parameter[0:207][7:0] ROM = {
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111100, // 2  *****
        8'b11000110, // 3 **   **
        8'b11000110, // 4 **   **
        8'b01100000, // 5  **
        8'b00111000, // 6   ***
        8'b00001100, // 7     **
        8'b00000110, // 8      **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b01111100, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

		  
        //E
		  8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2 *******
        8'b01100110, // 3  **  **
        8'b01100010, // 4  **   *
        8'b01101000, // 5  ** *
        8'b01111000, // 6  ****
        8'b01101000, // 7  ** *
        8'b01100000, // 8  **
        8'b01100010, // 9  **   *
        8'b01100110, // a  **  **
        8'b11111110, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
 
        //L
		  8'b00000000, // 0
        8'b00000000, // 1
        8'b11110000, // 2 ****
        8'b01100000, // 3  **
        8'b01100000, // 4  **
        8'b01100000, // 5  **
        8'b01100000, // 6  **
        8'b01100000, // 7  **
        8'b01100000, // 8  **
        8'b01100010, // 9  **   *
        8'b01100110, // a  **  **
        8'b11111110, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

		  //SPACE
	8'b00000000, // 0
	8'b00000000, // 1
	8'b00000000, // 2
	8'b00000000, // 3
	8'b00000000, // 4
	8'b00000000, // 5
	8'b00000000, // 6
	8'b00000000, // 7
	8'b00000000, // 8
	8'b00000000, // 9
	8'b00000000, // a
	8'b00000000, // b
	8'b00000000, // c
	8'b00000000, // d
	8'b00000000, // e
	8'b00000000, // f

        //M
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11000010, // 2 **    **
        8'b11100110, // 3 ***  ***
        8'b11111110, // 4 ********
        8'b11111110, // 5 ********
        8'b11011010, // 6 ** ** **
        8'b11000010, // 7 **    **
        8'b11000010, // 8 **    **
        8'b11000010, // 9 **    **
        8'b11000010, // a **    **
        8'b11000010, // b **    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

		  
		  
		  
        //O
		  8'b00000000, // 0
        8'b00000000, // 1
        8'b01111100, // 2  *****
        8'b11000110, // 3 **   **
        8'b11000110, // 4 **   **
        8'b11000110, // 5 **   **
        8'b11000110, // 6 **   **
        8'b11000110, // 7 **   **
        8'b11000110, // 8 **   **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b01111100, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

		  
		  
		 
        //D
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111000, // 2 *****
        8'b11000100, // 3 *   **
        8'b11000110, // 4 *   **
        8'b11000110, // 5 *   **
        8'b11000110, // 6 *   **
        8'b11000110, // 7 *   **
        8'b11000110, // 8 *   **
        8'b11000110, // 9 *   **
        8'b11000100, // a *   **
        8'b11111000, // b *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f	

		  
        //E
		  8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2 *******
        8'b01100110, // 3  **  **
        8'b01100010, // 4  **   *
        8'b01101000, // 5  ** *
        8'b01111000, // 6  ****
        8'b01101000, // 7  ** *
        8'b01100000, // 8  **
        8'b01100010, // 9  **   *
        8'b01100110, // a  **  **
        8'b11111110, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
		  
		  
		  
        //E
		  8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2 *******
        8'b01100110, // 3  **  **
        8'b01100010, // 4  **   *
        8'b01101000, // 5  ** *
        8'b01111000, // 6  ****
        8'b01101000, // 7  ** *
        8'b01100000, // 8  **
        8'b01100010, // 9  **   *
        8'b01100110, // a  **  **
        8'b11111110, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

		  //SPACE
	8'b00000000, // 0
	8'b00000000, // 1
	8'b00000000, // 2
	8'b00000000, // 3
	8'b00000000, // 4
	8'b00000000, // 5
	8'b00000000, // 6
	8'b00000000, // 7
	8'b00000000, // 8
	8'b00000000, // 9
	8'b00000000, // a
	8'b00000000, // b
	8'b00000000, // c
	8'b00000000, // d
	8'b00000000, // e
	8'b00000000, // f
		  
		  
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11000110, // 2 **   **
        8'b11100110, // 3 ***  **
        8'b11110110, // 4 **** **
        8'b11111110, // 5 *******
        8'b11011110, // 6 ** ****
        8'b11001110, // 7 **  ***
        8'b11000110, // 8 **   **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b11000110, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

		  
		  //SPACE
	8'b00000000, // 0
	8'b00000000, // 1
	8'b00000000, // 2
	8'b00000000, // 3
	8'b00000000, // 4
	8'b00000000, // 5
	8'b00000000, // 6
	8'b00000000, // 7
	8'b00000000, // 8
	8'b00000000, // 9
	8'b00000000, // a
	8'b00000000, // b
	8'b00000000, // c
	8'b00000000, // d
	8'b00000000, // e
	8'b00000000, // f
		 
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00010000, // 2    *
        8'b00111000, // 3   ***
        8'b01101100, // 4  ** **
        8'b11000110, // 5 **   **
        8'b11000110, // 6 **   **
        8'b11111110, // 7 *******
        8'b11000110, // 8 **   **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b11000110, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f	

		  
       

	};
	
	assign data = ROM[address];

endmodule 